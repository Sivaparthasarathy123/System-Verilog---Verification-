---------------OUTPUT----------------
Randomized Inputs: D = 1
 Generator Class 
Reset = 0| Input D = 1| output Q = 0
Randomized Inputs: D = 0
 Generator Class 
Reset = 1| Input D = 0| output Q = 0
Randomized Inputs: D = 0
 Generator Class 
Reset = 0| Input D = 0| output Q = 0
Randomized Inputs: D = 0
 Generator Class 
Reset = 1| Input D = 0| output Q = 0
Randomized Inputs: D = 1
 Generator Class 
Reset = 0| Input D = 1| output Q = 0
 Driver Class 
Reset = 0| Input D = 1| output Q = 0
 Monitor Class 
Reset = 0| Input D = 0| output Q = 0
PASS
 Scoreboard Class 
Reset = 0| Input D = 0| output Q = 0
 Driver Class 
Reset = 1| Input D = 0| output Q = 0
 Monitor Class 
Reset = 0| Input D = 1| output Q = 1
FAIL
 Scoreboard Class 
Reset = 0| Input D = 1| output Q = 1
 Driver Class 
Reset = 0| Input D = 0| output Q = 0
 Monitor Class 
Reset = 1| Input D = 0| output Q = 0
PASS
 Scoreboard Class 
Reset = 1| Input D = 0| output Q = 0
 Driver Class 
Reset = 1| Input D = 0| output Q = 0
 Monitor Class 
Reset = 0| Input D = 0| output Q = 0
PASS
 Scoreboard Class 
Reset = 0| Input D = 0| output Q = 0
 Driver Class 
Reset = 0| Input D = 1| output Q = 0
 Monitor Class 
Reset = 1| Input D = 0| output Q = 0
PASS
 Scoreboard Class 
Reset = 1| Input D = 0| output Q = 0
$finish at simulation time        60
