--- Generator Class ------
Time = 0 | Write Enable = 1 | Address = 0 | Data In = a9 | Data Out = 0
------ Monitor Class ------
Time = 5 | Write Enable = 0 | Address = 0 | Data In = 0 | Data Out = 0
[Scoreboard] PASS! Read 0 from Addr 0
------Scoreboard Class---
---
Time = 5 | Write Enable = 0 | Address = 0 | Data In = 0 | Data Out = 0
---
--- Generator Class ------
Time = 5 | Write Enable = 1 | Address = 7 | Data In = b8 | Data Out = 0
------ Driver Class ------
Time = 10 | Write Enable = 1 | Address = 0 | Data In = a9 | Data Out = 0
------ Monitor Class ------
Time = 15 | Write Enable = 1 | Address = 0 | Data In = a9 | Data Out = 0
[Scoreboard] Model Write a9 to Addr 0
[Scoreboard] PASS! Read 0 from Addr 0
------Scoreboard Class---
---
Time = 15 | Write Enable = 1 | Address = 0 | Data In = a9 | Data Out = 0
---
--- Generator Class ------
Time = 15 | Write Enable = 1 | Address = 0 | Data In = ee | Data Out = 0
------ Driver Class ------
Time = 20 | Write Enable = 1 | Address = 7 | Data In = b8 | Data Out = 0
------ Monitor Class ------
Time = 25 | Write Enable = 1 | Address = 7 | Data In = b8 | Data Out = 0
[Scoreboard] Model Write b8 to Addr 7
[Scoreboard] PASS! Read 0 from Addr 7
------Scoreboard Class---
---
Time = 25 | Write Enable = 1 | Address = 7 | Data In = b8 | Data Out = 0
---
--- Generator Class ------
Time = 25 | Write Enable = 1 | Address = 1 | Data In = aa | Data Out = 0
------ Driver Class ------
Time = 30 | Write Enable = 1 | Address = 0 | Data In = ee | Data Out = 0
------ Monitor Class ------
Time = 35 | Write Enable = 1 | Address = 0 | Data In = ee | Data Out = a9
[Scoreboard] Model Write ee to Addr 0
[Scoreboard] PASS! Read a9 from Addr 0
------Scoreboard Class---
---
Time = 35 | Write Enable = 1 | Address = 0 | Data In = ee | Data Out = a9
---
--- Generator Class ------
Time = 35 | Write Enable = 1 | Address = 4 | Data In = ab | Data Out = 0
------ Driver Class ------
Time = 40 | Write Enable = 1 | Address = 1 | Data In = aa | Data Out = 0
------ Monitor Class ------
Time = 45 | Write Enable = 1 | Address = 1 | Data In = aa | Data Out = 0
[Scoreboard] Model Write aa to Addr 1
[Scoreboard] PASS! Read 0 from Addr 1
------Scoreboard Class---
---
Time = 45 | Write Enable = 1 | Address = 1 | Data In = aa | Data Out = 0
---
--- Generator Class ------
Time = 45 | Write Enable = 1 | Address = 2 | Data In = b4 | Data Out = 0
------ Driver Class ------
Time = 50 | Write Enable = 1 | Address = 4 | Data In = ab | Data Out = 0
------ Monitor Class ------
Time = 55 | Write Enable = 1 | Address = 4 | Data In = ab | Data Out = 0
[Scoreboard] Model Write ab to Addr 4
[Scoreboard] PASS! Read 0 from Addr 4
------Scoreboard Class---
---
Time = 55 | Write Enable = 1 | Address = 4 | Data In = ab | Data Out = 0
---
--- Generator Class ------
Time = 55 | Write Enable = 1 | Address = 7 | Data In = f9 | Data Out = 0
------ Driver Class ------
Time = 60 | Write Enable = 1 | Address = 2 | Data In = b4 | Data Out = 0
------ Monitor Class ------
Time = 65 | Write Enable = 1 | Address = 2 | Data In = b4 | Data Out = 0
[Scoreboard] Model Write b4 to Addr 2
[Scoreboard] PASS! Read 0 from Addr 2
------Scoreboard Class---
---
Time = 65 | Write Enable = 1 | Address = 2 | Data In = b4 | Data Out = 0
---
--- Generator Class ------
Time = 65 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 0
------ Driver Class ------
Time = 70 | Write Enable = 1 | Address = 7 | Data In = f9 | Data Out = 0
------ Monitor Class ------
Time = 75 | Write Enable = 1 | Address = 7 | Data In = f9 | Data Out = b8
[Scoreboard] Model Write f9 to Addr 7
[Scoreboard] PASS! Read b8 from Addr 7
------Scoreboard Class---
---
Time = 75 | Write Enable = 1 | Address = 7 | Data In = f9 | Data Out = b8
---
--- Generator Class ------
Time = 75 | Write Enable = 1 | Address = 2 | Data In = f6 | Data Out = 0
------ Driver Class ------
Time = 80 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 0
------ Monitor Class ------
Time = 85 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = aa
[Scoreboard] Model Write 1f to Addr 1
[Scoreboard] PASS! Read aa from Addr 1
------Scoreboard Class---
---
Time = 85 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = aa
---
--- Generator Class ------
Time = 85 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 0
------ Driver Class ------
Time = 90 | Write Enable = 1 | Address = 2 | Data In = f6 | Data Out = 0
------ Monitor Class ------
Time = 95 | Write Enable = 1 | Address = 2 | Data In = f6 | Data Out = b4
[Scoreboard] Model Write f6 to Addr 2
[Scoreboard] PASS! Read b4 from Addr 2
------Scoreboard Class---
---
Time = 95 | Write Enable = 1 | Address = 2 | Data In = f6 | Data Out = b4
---
--- Generator Class ------
Time = 95 | Write Enable = 1 | Address = 2 | Data In = f5 | Data Out = 0
------ Driver Class ------
Time = 100 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 0
------ Monitor Class ------
Time = 105 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 1f
[Scoreboard] Model Write 1f to Addr 1
[Scoreboard] PASS! Read 1f from Addr 1
------Scoreboard Class---
---
Time = 105 | Write Enable = 1 | Address = 1 | Data In = 1f | Data Out = 1f
---
--- Generator Class ------
Time = 105 | Write Enable = 1 | Address = 6 | Data In = 55 | Data Out = 0
------ Driver Class ------
Time = 110 | Write Enable = 1 | Address = 2 | Data In = f5 | Data Out = 0
------ Monitor Class ------
Time = 115 | Write Enable = 1 | Address = 2 | Data In = f5 | Data Out = f6
[Scoreboard] Model Write f5 to Addr 2
[Scoreboard] PASS! Read f6 from Addr 2
------Scoreboard Class---
---
Time = 115 | Write Enable = 1 | Address = 2 | Data In = f5 | Data Out = f6
---
--- Generator Class ------
Time = 115 | Write Enable = 1 | Address = 5 | Data In = 2b | Data Out = 0
------ Driver Class ------
Time = 120 | Write Enable = 1 | Address = 6 | Data In = 55 | Data Out = 0
------ Monitor Class ------
Time = 125 | Write Enable = 1 | Address = 6 | Data In = 55 | Data Out = 0
[Scoreboard] Model Write 55 to Addr 6
[Scoreboard] PASS! Read 0 from Addr 6
------Scoreboard Class---
---
Time = 125 | Write Enable = 1 | Address = 6 | Data In = 55 | Data Out = 0
---
--- Generator Class ------
Time = 125 | Write Enable = 1 | Address = 6 | Data In = 13 | Data Out = 0
------ Driver Class ------
Time = 130 | Write Enable = 1 | Address = 5 | Data In = 2b | Data Out = 0
------ Monitor Class ------
Time = 135 | Write Enable = 1 | Address = 5 | Data In = 2b | Data Out = 0
[Scoreboard] Model Write 2b to Addr 5
[Scoreboard] PASS! Read 0 from Addr 5
------Scoreboard Class---
---
Time = 135 | Write Enable = 1 | Address = 5 | Data In = 2b | Data Out = 0
---
--- Generator Class ------
Time = 135 | Write Enable = 1 | Address = 1 | Data In = 7d | Data Out = 0
------ Driver Class ------
Time = 140 | Write Enable = 1 | Address = 6 | Data In = 13 | Data Out = 0
------ Monitor Class ------
Time = 145 | Write Enable = 1 | Address = 6 | Data In = 13 | Data Out = 55
[Scoreboard] Model Write 13 to Addr 6
[Scoreboard] PASS! Read 55 from Addr 6
------Scoreboard Class---
---
Time = 145 | Write Enable = 1 | Address = 6 | Data In = 13 | Data Out = 55
------ Driver Class ------
Time = 150 | Write Enable = 1 | Address = 1 | Data In = 7d | Data Out = 0
--- Final Verification Success ---
$finish called from file "test.sv", line 12.
$finish at simulation time                  170
