Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Dec 29 10:48 2025
Passed value: a=0 b=0 cin=0 sum=0 carry=0
Passed value: a=1 b=1 cin=1 sum=1 carry=1
Passed value: a=1 b=0 cin=1 sum=0 carry=1
$finish at simulation time               
