Randomized Inputs: Reset = 0| Enable = 1
Generator Class
Time = 0| Reset = 0| Enable = 1| Output Q = 0
Randomized Inputs: Reset = 1| Enable = 0
Generator Class
Time = 5| Reset = 1| Enable = 0| Output Q = 0
Driver Class
Time = 5| Reset = 0| Enable = 1| Output Q = 0
Monitor Class
Time = 5| Reset = 0| Enable = 1| Output Q = 1
PASS: Expected Output Q = 1| Output Q = 1
Randomized Inputs: Reset = 0| Enable = 0
Generator Class
Time = 10| Reset = 0| Enable = 0| Output Q = 0
Randomized Inputs: Reset = 1| Enable = 0
Generator Class
Time = 15| Reset = 1| Enable = 0| Output Q = 0
Driver Class
Time = 15| Reset = 1| Enable = 0| Output Q = 0
Monitor Class
Time = 15| Reset = 0| Enable = 0| Output Q = 6
PASS: Expected Output Q = 6| Output Q = 6
Randomized Inputs: Reset = 0| Enable = 1
Generator Class
Time = 20| Reset = 0| Enable = 1| Output Q = 0
Driver Class
Time = 25| Reset = 0| Enable = 0| Output Q = 0
Monitor Class
Time = 25| Reset = 0| Enable = 0| Output Q = 6
PASS: Expected Output Q = 6| Output Q = 6
Driver Class
Time = 35| Reset = 1| Enable = 0| Output Q = 0
Monitor Class
Time = 35| Reset = 1| Enable = 0| Output Q = 0
PASS: Expected Output Q = 0| Output Q = 0
Driver Class
Time = 45| Reset = 0| Enable = 1| Output Q = 0
Monitor Class
Time = 45| Reset = 0| Enable = 1| Output Q = 1
PASS: Expected Output Q = 1| Output Q = 1
$finish at simulation time                   55
