--------------- Output -------------------
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 169 (10101001) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 184 (10111000) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 238 (11101110) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 170 (10101010) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 171 (10101011) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 180 (10110100) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 249 (11111001) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 31 (11111) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 246 (11110110) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: w_rst = 0 | w_en = 1
----  Generator class for Write Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 31 (11111) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
Time = 0 | Randomized Inputs: r_rst = 0 | r_en = 1
----  Generator class for Read Operation  ----
Time = 0 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Write Value to Driver  ----
Time = 5000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 169 (10101001) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 5000 | w_rst = 1 | r_rst = 0 | w_en = 0 | r_en = 0 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_RESET] Time=5000 | Queue Cleared
----  Write Value to Driver  ----
Time = 15000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 184 (10111000) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 15000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 169 (10101001) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_WRITE] Time=15000 | Data In: 169
----  Write Value to Driver  ----
Time = 25000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 238 (11101110) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 25000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 184 (10111000) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_WRITE] Time=25000 | Data In: 184
----  Write Value to Driver  ----
Time = 35000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 170 (10101010) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 35000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 238 (11101110) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_WRITE] Time=35000 | Data In: 238
----  Write Value to Driver  ----
Time = 45000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 171 (10101011) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 45000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 170 (10101010) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_WRITE] Time=45000 | Data In: 170
----  Write Value to Driver  ----
Time = 55000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 180 (10110100) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 55000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 171 (10101011) | Data out = 0 (0) | Full = 0 | Empty = 0
[SCB_WRITE] Time=55000 | Data In: 171
----  Write Value to Driver  ----
Time = 65000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 249 (11111001) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 65000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 180 (10110100) | Data out = 0 (0) | Full = 1 | Empty = 0
----  Write Value to Driver  ----
Time = 75000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 31 (11111) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 75000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 249 (11111001) | Data out = 0 (0) | Full = 1 | Empty = 0
----  Write Value to Driver  ----
Time = 85000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 246 (11110110) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 85000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 31 (11111) | Data out = 0 (0) | Full = 1 | Empty = 0
----  Write Value to Driver  ----
Time = 95000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 31 (11111) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 95000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 0 | Data in = 246 (11110110) | Data out = 0 (0) | Full = 1 | Empty = 0
----   Read Value to Driver  ----
Time = 105000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 105000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 0 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----   Read Value to Driver  ----
Time = 115000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 115000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 169 (10101001) | Full = 0 | Empty = 0
[SCB_PASS] Got: 169
----   Read Value to Driver  ----
Time = 125000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 125000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 184 (10111000) | Full = 0 | Empty = 0
[SCB_PASS] Got: 184
----   Read Value to Driver  ----
Time = 135000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 135000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 238 (11101110) | Full = 0 | Empty = 0
[SCB_PASS] Got: 238
----   Read Value to Driver  ----
Time = 145000 | w_rst = 0 | r_rst = 0 | w_en = 1 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 145000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 170 (10101010) | Full = 0 | Empty = 0
[SCB_PASS] Got: 170
----   Read Value to Driver  ----
Time = 155000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 155000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 171 (10101011) | Full = 0 | Empty = 0
[SCB_PASS] Got: 171
----   Read Value to Driver  ----
Time = 165000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 165000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 180 (10110100) | Full = 0 | Empty = 0
----   Read Value to Driver  ----
Time = 175000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 175000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 31 (11111) | Full = 0 | Empty = 0
----   Read Value to Driver  ----
Time = 185000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 185000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----   Read Value to Driver  ----
Time = 195000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
----  Value to Monitor  ----
Time = 195000 | w_rst = 0 | r_rst = 0 | w_en = 0 | r_en = 1 | Data in = 0 (0) | Data out = 0 (0) | Full = 0 | Empty = 0
$finish called from file "testbench.sv", line 44.
$finish at simulation time              1020000
