// Interface creation
interface f_adder;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic carry;
  
endinterface
